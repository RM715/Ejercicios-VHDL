----------------------------------------------------------------------------------
-- Company: 
-- Engineer: 
-- 
-- Create Date:    22:37:29 05/18/2022 
-- Design Name: 
-- Module Name:    Promedio2 - Behavioral 
-- Project Name: 
-- Target Devices: 
-- Tool versions: 
-- Description: 
--
-- Dependencies: 
--
-- Revision: 
-- Revision 0.01 - File Created
-- Additional Comments: 
--
----------------------------------------------------------------------------------
library IEEE;
use IEEE.STD_LOGIC_1164.ALL;

-- Uncomment the following library declaration if using
-- arithmetic functions with Signed or Unsigned values
--use IEEE.NUMERIC_STD.ALL;

-- Uncomment the following library declaration if instantiating
-- any Xilinx primitives in this code.
--library UNISIM;
--use UNISIM.VComponents.all;

entity Promedio2 is
    Port ( A : in  STD_LOGIC_VECTOR (0 to 3);
           B : in  STD_LOGIC_VECTOR (0 to 3);
           C : out  STD_LOGIC_VECTOR (0 to 3));
end Promedio2;

architecture Behavioral of Promedio2 is

begin


end Behavioral;

